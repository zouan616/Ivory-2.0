Buck_Converter.cir

.MODEL SWI SW(VT=4.5V VH=0V RON=0.0001 ROFF=1MEG)
.MODEL DSCH D(IS=0.0002 RS=0.0001 CJO=5e-10)

*SWITCH DRIVER 
VCTRL1 101 0 PULSE(-5V 5V 0.00NS 0NS 0NS 2NS 0.004US)
VCTRL2 102 0 PULSE(-5V 5V 0.125NS 0NS 0NS 2NS 0.004US)
VCTRL3 103 0 PULSE(-5V 5V 0.250NS 0NS 0NS 2NS 0.004US)
VCTRL4 104 0 PULSE(-5V 5V 0.375NS 0NS 0NS 2NS 0.004US)
VCTRL5 105 0 PULSE(-5V 5V 0.500NS 0NS 0NS 2NS 0.004US)
VCTRL6 106 0 PULSE(-5V 5V 0.625NS 0NS 0NS 2NS 0.004US)
VCTRL7 107 0 PULSE(-5V 5V 0.750NS 0NS 0NS 2NS 0.004US)
VCTRL8 108 0 PULSE(-5V 5V 0.875NS 0NS 0NS 2NS 0.004US)
VCTRL9 109 0 PULSE(-5V 5V 1.00NS 0NS 0NS 2US 0.004US)
VCTRL10 110 0 PULSE(-5V 5V 1.125NS 0NS 0NS 2NS 0.004US)
VCTRL11 111 0 PULSE(-5V 5V 1.250NS 0NS 0NS 2NS 0.004US)
VCTRL12 112 0 PULSE(-5V 5V 1.375NS 0NS 0NS 2NS 0.004US)
VCTRL13 113 0 PULSE(-5V 5V 1.500NS 0NS 0NS 2NS 0.004US)
VCTRL14 114 0 PULSE(-5V 5V 1.625NS 0NS 0NS 2NS 0.004US)
VCTRL15 115 0 PULSE(-5V 5V 1.750NS 0NS 0NS 2NS 0.004US)
VCTRL16 116 0 PULSE(-5V 5V 1.875NS 0NS 0NS 2NS 0.004US)


*INPUT VOLTAGE
VIN 1 0 SIN(0 1 1000000000 0ns 0 0)

* CONVERTER 1
SW1 1 2	101 0 SWI
SW1b2 0 2 0 101 SWI
L1 2 3 0.011uH
* CONVERTER 2
SW2 1 4	102 0 SWI
SW2b2 0 4 0 102 SWI
L2 4 3 0.011uH
* CONVERTER 3
SW3 1 5	103 0 SWI
SW3b2 0 5 0 103 SWI
L3 5 3 0.011uH
* CONVERTER 4
SW4 1 6	104 0 SWI
SW4b2 0 6 0 104 SWI
L4 6 3 0.011uH
* CONVERTER 5
SW5 1 7	105 0 SWI
SW5b2 0 7 0 105 SWI
L5 7 3 0.011uH
* CONVERTER 6
SW6 1 8	106 0 SWI
SW6b2 0 8 0 106 SWI
L6 8 3 0.011uH
* CONVERTER 7
SW7 1 9	107 0 SWI
SW7b2 0 9 0 107 SWI
L7 9 3 0.011uH
* CONVERTER 8
SW8 1 10 108 0 SWI
SW8b2 0 10 0 108 SWI
L8 10 3 0.011uH
* CONVERTER 9
SW9 1 11 109 0 SWI
SW9b2 0 11 0 109 SWI
L9 11 3 0.011uH
* CONVERTER 10
SW10 1 12 110 0 SWI
SW10b2 0 12 0 110 SWI
L10 12 3 0.011uH
* CONVERTER 11
SW11 1 13 111 0 SWI
SW11b2 0 13 0 111 SWI
L11 13 3 0.011uH
* CONVERTER 12
SW12 1 14 112 0 SWI
SW12b2 0 14 0 112 SWI
L12 14 3 0.011uH
* CONVERTER 13
SW13 1 15 113 0 SWI
SW13b2 0 15 0 113 SWI
L13 15 3 0.011uH
* CONVERTER 14
SW14 1 16 114 0 SWI
SW14b2 0 16 0 114 SWI
L14 16 3 0.011uH
* CONVERTER 15
SW15 1 17 115 0 SWI
SW15b2 0 17 0 115 SWI
L15 17 3 0.011uH
* CONVERTER 16
SW16 1 18 116 0 SWI
SW16b2 0 18 0 116 SWI
L16 18 3 0.011uH




C1 3 0 0.096UF

*LOAD
RL 3 0 5

.TRAN 0.0001US 10US

.END

