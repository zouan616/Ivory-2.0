Buck_Converter_8.cir

.MODEL SWI SW(VT=4.5V VH=0V RON=0.0001 ROFF=1MEG)
.MODEL DSCH D(IS=0.0002 RS=0.0001 CJO=5e-10)

*SWITCH DRIVER 
VCTRL1 101 0 PULSE(-5V 5V 0.00125US 0NS 0NS 0.005US 0.01US)
VCTRL2 102 0 PULSE(-5V 5V 0.0025 0NS 0NS 0.005US 0.01US)
VCTRL3 103 0 PULSE(-5V 5V 0.00375US 0NS 0NS 0.005US 0.01US)
VCTRL4 104 0 PULSE(-5V 5V 0.005US 0NS 0NS 0.005US 0.01US)
VCTRL5 105 0 PULSE(-5V 5V 0.00625NS 0NS 0NS 0.005US 0.01US)
VCTRL6 106 0 PULSE(-5V 5V 0.0075US 0NS 0NS 0.005US 0.01US)
VCTRL7 107 0 PULSE(-5V 5V 0.00875US 0NS 0NS 0.005US 0.01US)
VCTRL8 108 0 PULSE(-5V 5V 0.01US 0NS 0NS 0.005US 0.01US)



*INPUT VOLTAGE
VIN 1 0 SIN(0 1 7000000 0ns 0 0)

* CONVERTER 1
SW1 1 2	101 0 SWI
SW1b2 0 2 0 101 SWI
L1 2 3 1.8nH
* CONVERTER 2
SW2 1 4	102 0 SWI
SW2b2 0 4 0 102 SWI
L2 4 3 1.8nH
* CONVERTER 3
SW3 1 5	103 0 SWI
SW3b2 0 5 0 103 SWI
L3 5 3 1.8nH
* CONVERTER 4
SW4 1 6	104 0 SWI
SW4b2 0 6 0 104 SWI
L4 6 3 1.8nH
* CONVERTER 5
SW5 1 7	105 0 SWI
SW5b2 0 7 0 105 SWI
L5 7 3 1.8nH
* CONVERTER 6
SW6 1 8	106 0 SWI
SW6b2 0 8 0 106 SWI
L6 8 3 1.8nH
* CONVERTER 7
SW7 1 9	107 0 SWI
SW7b2 0 9 0 107 SWI
L7 9 3 1.8nH
* CONVERTER 8
SW8 1 10 108 0 SWI
SW8b2 0 10 0 108 SWI
L8 10 3 1.8nH





C1 3 0 8.8UF

*LOAD
RL 3 0 1

.TRAN 0.0001US 100US

.END

