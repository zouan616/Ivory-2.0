Buck_Converter.cir

.MODEL SWI SW(VT=4.5V VH=0V RON=0.0001 ROFF=1MEG)
.MODEL DSCH D(IS=0.0002 RS=0.0001 CJO=5e-10)

*SWITCH DRIVER 
VCTRL1 101 0 PULSE(0V 5V 1NS 1NS 1NS 0.2US 2US)
VCTRL2 102 0 PULSE(0V 5V 0.125US 1NS 1NS 0.2US 2US)
VCTRL3 103 0 PULSE(0V 5V 0.25US 1NS 1NS 0.2US 2US)
VCTRL4 104 0 PULSE(0V 5V 0.375US 1NS 1NS 0.2US 2US)
VCTRL5 105 0 PULSE(0V 5V 0.50US 1NS 1NS 0.2US 2US)
VCTRL6 106 0 PULSE(0V 5V 0.625US 1NS 1NS 0.2US 2US)
VCTRL7 107 0 PULSE(0V 5V 0.75US 1NS 1NS 0.2US 2US)
VCTRL8 108 0 PULSE(0V 5V 0.875US 1NS 1NS 0.2US 2US)
VCTRL9 109 0 PULSE(0V 5V 1.000US 1NS 1NS 0.2US 2US)
VCTRL10 110 0 PULSE(0V 5V 1.125US 1NS 1NS 0.2US 2US)
VCTRL11 111 0 PULSE(0V 5V 1.25US 1NS 1NS 0.2US 2US)
VCTRL12 112 0 PULSE(0V 5V 1.375US 1NS 1NS 0.2US 2US)
VCTRL13 113 0 PULSE(0V 5V 1.50US 1NS 1NS 0.2US 2US)
VCTRL14 114 0 PULSE(0V 5V 1.625US 1NS 1NS 0.2US 2US)
VCTRL15 115 0 PULSE(0V 5V 1.750US 1NS 1NS 0.2US 2US)
VCTRL16 116 0 PULSE(0V 5V 1.875USS 1NS 1NS 0.2US 2US)


*INPUT VOLTAGE
VIN 1 0 SIN(0 1 1000 1ns 0 0)

* CONVERTER 1
SW1 1 2	101 0 SWI
D1 0 2 DSCH
L1 2 3 0.1mH
* CONVERTER 2
SW2 1 4	102 0 SWI
D2 0 4 DSCH
L2 4 3 0.1mH
* CONVERTER 3
SW3 1 5	103 0 SWI
D3 0 5 DSCH
L3 5 3 0.1mH
* CONVERTER 4
SW4 1 6	104 0 SWI
D4 0 6 DSCH
L4 6 3 0.1mH
* CONVERTER 5
SW5 1 7	105 0 SWI
D5 0 7 DSCH
L5 7 3 0.1mH
* CONVERTER 6
SW6 1 8	106 0 SWI
D6 0 8 DSCH
L6 8 3 0.1mH
* CONVERTER 7
SW7 1 9	107 0 SWI
D7 0 9 DSCH
L7 9 3 0.1mH
* CONVERTER 8
SW8 1 10 108 0 SWI
D8 0 10 DSCH
L8 10 3 0.1mH
* CONVERTER 9
SW9 1 11 109 0 SWI
D9 0 11 DSCH
L9 11 3 0.1mH
* CONVERTER 10
SW10 1 12 110 0 SWI
D10 0 12 DSCH
L10 12 3 0.1mH
* CONVERTER 11
SW11 1 13 111 0 SWI
D11 0 13 DSCH
L11 13 3 0.1mH
* CONVERTER 12
SW12 1 14 112 0 SWI
D12 0 14 DSCH
L12 14 3 0.1mH
* CONVERTER 13
SW13 1 15 113 0 SWI
D13 0 15 DSCH
L13 15 3 0.1mH
* CONVERTER 14
SW14 1 16 114 0 SWI
D14 0 16 DSCH
L14 16 3 0.1mH
* CONVERTER 15
SW15 1 17 115 0 SWI
D15 0 17 DSCH
L15 17 3 0.1mH
* CONVERTER 16
SW16 1 18 116 0 SWI
D16 0 18 DSCH
L16 18 3 0.1mH




C1 3 0 0.10UF

*LOAD
RL 3 0 1

.TRAN 0.0001US 5000US

.END

