Buck_Converter_6.cir

.MODEL SWI SW(VT=4.5V VH=0V RON=0.01 ROFF=1MEG)
.MODEL DSCH D(IS=0.0002 RS=0.01 CJO=5e-10)

*SWITCH DRIVER 
VCTRL1 101 0 PULSE(0V 5V 1NS 1NS 1NS 1US 2US)
VCTRL2 102 0 PULSE(0V 5V 0.4US 1NS 1NS 1US 2US)
VCTRL3 103 0 PULSE(0V 5V 0.8US 1NS 1NS 1US 2US)
VCTRL4 104 0 PULSE(0V 5V 1.2US 1NS 1NS 1US 2US)
VCTRL5 105 0 PULSE(0V 5V 1.6US 1NS 1NS 1US 2US)
VCTRL6 106 0 PULSE(0V 5V 1.6US 1NS 1NS 1US 2US)

*INPUT VOLTAGE
VIN 1 0 SIN(10 1 500000 1ns 0 0)

* CONVERTER 1
SW1 1 2	101 0 SWI
D1 0 2 DSCH
L1 2 3 0.05mH
* CONVERTER 2
SW2 1 4	102 0 SWI
D2 0 4 DSCH
L2 4 3 0.02mH
* CONVERTER 3
SW3 1 5	103 0 SWI
D3 0 5 DSCH
L3 5 3 0.02mH
* CONVERTER 4
SW4 1 6	104 0 SWI
D4 0 6 DSCH
L4 6 3 0.02mH
SW5 1 7	105 0 SWI
D5 0 7 DSCH
L5 7 3 0.02mH
SW6 1 8	106 0 SWI
D6 0 8 DSCH
L6 8 3 0.02mH


C1 3 0 0.10UF

*LOAD
RL 3 0 1

.TRAN 0.0001US 1000US

.END

