Buck_Converter.cir

.MODEL SWI SW(VT=4.5V VH=0V RON=0.01 ROFF=1MEG)
.MODEL DSCH D(IS=0.0002 RS=0.01 CJO=5e-10)

*SWITCH DRIVER 
VCTRL 10 0 PULSE(0V 5V 1NS 1NS 1NS 1US 2US)


*INPUT VOLTAGE
VIN 1 0 SIN(10 1 100000 1ns 0 0)

* CONVERTER
SW1 1 2	10 0 SWI
D1 0 2 DSCH
L1 2 3 0.1mH
C1 3 0 0.10UF

*LOAD
RL 3 0 1

.TRAN 0.01US 100000US

.END
