Buck_Converter_2.cir

.MODEL SWI SW(VT=4.5V VH=0V RON=0.01 ROFF=1MEG)
.MODEL DSCH D(IS=0.0002 RS=0.01 CJO=5e-10)

*SWITCH DRIVER 
VCTRL1 10 0 PULSE(0V 5V 1NS 1NS 1NS 0.2US 2US)
VCTRL2 11 0 PULSE(0V 5V 1US 1NS 1NS 0.2US 2US)


*INPUT VOLTAGE
VIN 1 0 SIN(10 1 500000 1ns 0 0)

* CONVERTER phase 1
SW1 1 2	10 0 SWI
D1 0 2 DSCH
L1 2 3 0.05mH
* CONVERTER phase 2
SW2 1 4	11 0 SWI
D2 0 4 DSCH
L2 4 3 0.05mH



C1 3 0 0.10UF

*LOAD
RL 3 0 1

.TRAN 0.0001US 2000US

.END
