Buck_Converter_1_model.cir

.MODEL SWI SW(VT=4.5V VH=0V RON=1e-8 ROFF=1MEG)
.MODEL DSCH D(IS=0.0002 RS=1e-8 CJO=5e-10)

*SWITCH DRIVER 
VCTRL1 101 0 PULSE(0V 5V 1NS 1NS 1NS 0.01US 0.01US)



*INPUT VOLTAGE
*VIN 1 0 PULSE(10 1 10us 1ns 1ns 1 2 0)
VIN 1 0 DC 1.1

* CONVERTER 1
SW1 1 2	101 0 SWI
D1 0 2 DSCH
L1 2 3 0.1uH





C1 3 0 0.5UF

*LOAD
RL 3 0 0.5

.TRAN 0.0001US 100US

.END

