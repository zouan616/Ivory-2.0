Buck_Converter_4.cir

.MODEL SWI SW(VT=4.5V VH=0V RON=0.001 ROFF=1MEG)
.MODEL DSCH D(IS=0.0002 RS=0.001 CJO=5e-10)

*SWITCH DRIVER 
VCTRL1 101 0 PULSE(0V 5V 1NS 1NS 1NS 0.2US 2US)
VCTRL2 102 0 PULSE(0V 5V 0.5US 1NS 1NS 0.2US 2US)
VCTRL3 103 0 PULSE(0V 5V 1.0US 1NS 1NS 0.2US 2US)
VCTRL4 104 0 PULSE(0V 5V 1.5US 1NS 1NS 0.2US 2US)



*INPUT VOLTAGE
VIN 1 0 SIN(10 1 50000000 1ns 0 0)

* CONVERTER 1
SW1 1 2	101 0 SWI
D1 0 2 DSCH
L1 2 3 0.1mH
* CONVERTER 2
SW2 1 4	102 0 SWI
D2 0 4 DSCH
L2 4 3 0.1mH
* CONVERTER 3
SW3 1 5	103 0 SWI
D3 0 5 DSCH
L3 5 3 0.1mH
* CONVERTER 4
SW4 1 6	104 0 SWI
D4 0 6 DSCH
L4 6 3 0.1mH



C1 3 0 0.10UF

*LOAD
RL 3 0 1

.TRAN 0.001US 2000US

.END

