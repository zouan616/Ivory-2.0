Buck_Converter_10.cir

.MODEL SWI SW(VT=4.5V VH=0V RON=1e-7 ROFF=1MEG)
.MODEL DSCH D(IS=0.0002 RS=1e-7 CJO=5e-11)

*SWITCH DRIVER 
VCTRL1 101 0 PULSE(0V 5V 0NS 1NS 1NS 0.01US 0.05US)
VCTRL2 102 0 PULSE(0V 5V 0.005US 1NS 1NS 0.01US 0.05US)
VCTRL3 103 0 PULSE(0V 5V 0.01US 1NS 1NS 0.01US 0.05US)
VCTRL4 104 0 PULSE(0V 5V 0.015US 1NS 1NS 0.01US 0.05US)
VCTRL5 105 0 PULSE(0V 5V 0.02US 1NS 1NS 0.01US 0.05US)
VCTRL6 106 0 PULSE(0V 5V 0.025US 1NS 1NS 0.01US 0.05US)
VCTRL7 107 0 PULSE(0V 5V 0.03US 1NS 1NS 0.01US 0.05US)
VCTRL8 108 0 PULSE(0V 5V 0.035US 1NS 1NS 0.01US 0.05US)
VCTRL9 109 0 PULSE(0V 5V 0.04US 1NS 1NS 0.01US 0.05US)
VCTRL10 110 0 PULSE(0V 5V 0.045US 1NS 1NS 0.01US 0.05US)

*INPUT VOLTAGE
VIN 1 0 DC 5.42

* CONVERTER 1
SW1 1 2	101 0 SWI
D1 0 2 DSCH
L1 2 3 1uH
* CONVERTER 2
SW2 1 4	102 0 SWI
D2 0 4 DSCH
L2 4 3 1uH
* CONVERTER 3
SW3 1 5	103 0 SWI
D3 0 5 DSCH
L3 5 3 1uH
* CONVERTER 4
SW4 1 6	104 0 SWI
D4 0 6 DSCH
L4 6 3 1uH
* CONVERTER 5
SW5 1 7	105 0 SWI
D5 0 7 DSCH
L5 7 3 1uH
* CONVERTER 6
SW6 1 8	106 0 SWI
D6 0 8 DSCH
L6 8 3 1uH
* CONVERTER 7
SW7 1 9	107 0 SWI
D7 0 9 DSCH
L7 9 3 1uH
* CONVERTER 8
SW8 1 10 108 0 SWI
D8 0 10 DSCH
L8 10 3 1uH
* CONVERTER 9
SW9 1 11 109 0 SWI
D9 0 11 DSCH
L9 11 3 1uH
* CONVERTER 10
SW10 1 12 110 0 SWI
D10 0 12 DSCH
L10 12 3 1uH


C1 3 0 0.5UF

*LOAD
RL 3 0 0.5

.TRAN 0.0001US 100US

.END

